Full Rectifier

* .model <model name> D (N = 1m, Is = 1nA)
.MODEL 1N4148  D(Is=0.1p Rs=1.6 CJO=2p Tt=12n Bv=100 Ibv=0.1p)

Vin 3 2 SIN(0, 5, 1)
D1 3 1 1N4148
D2 0 2 1N4148
D3 0 3 1N4148
D4 2 1 1N4148
R1 1 0 1K

* .DC lin Vin -5 5 0.01
.tran 0.01 3

.end
