Simple Diode Circuit

* .model <model name> D (N = 1m, Is = 1nA)
.MODEL 1N4148  D(Is=0.1p Rs=1.6 CJO=2p Tt=12n Bv=100 Ibv=0.1p)

*Vin 1 0 SIN(0, 5, 1)
*R1 2 0 1k
*D1 1 2 1N4148

Vin 1 0 DC 5V
V1 3 0 DC 2
R1 3 2 1k
D1 2 1 1N4148

.DC lin Vin 0 5 0.01
* .tran 0.01 3 0

.end
