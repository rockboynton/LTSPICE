Full-wave rectifier and filter capacitor stages of a power supply

* accepts a 5V peak transformed secondary voltage V2 and limits the ripple
* voltage to 5% if RL = 2K

.MODEL 1N4148  D(Is=0.1p Rs=1.6 CJO=2p Tt=12n Bv=100 Ibv=0.1p)

Vin 1 3 SIN(0, 5, 60)
D1 1 2 1N4148
D2 0 3 1N4148
D3 0 1 1N4148
D4 3 2 1N4148
C1 2 0 83.33uF
R1 2 0 2k

.tran 1us 100ms

.end
