Lab rectifier

.MODEL 1N4148  D(Is=0.1p Rs=1.6 CJO=2p Tt=12n Bv=100 Ibv=0.1p)

V1 1 0 1
D1 1 2 1N4148
D2 3 2 1N4148
R1 2 0 2k
E2 0 3 1 0 1

.dc V1 -5 5 1

.end
